創世神
Priest
96
100
1
0
1
2
back:
staff
backend
