﻿你好
Priest
100
100
1
0
1
87
back:
staff
backend
staff
none
none
none
