小可愛
Swordsman
100
100
1
10
2
900032
back:
GodSword
backend
